`timescale 1ns / 1ps	//!< <time unit> / <time precision>

`include "TD4.v"

module TD4_testbench();

endmodule